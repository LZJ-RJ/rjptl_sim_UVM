`timescale 1ps/1ps
package rjptl_pkg_dut;

// Part 1 - Official UVM
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "enum_dut.svh"

endpackage