// Sequence
`include "super_like_rj_seq.sv"

// Test
`include "base_test.sv"
`include "super_like_rj_test_case.sv"