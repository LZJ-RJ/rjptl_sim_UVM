class super_like_rj_seq extends rj_sequence;
    `uvm_object_utils(super_like_rj_seq)
    function new(string name = "super_like_rj_seq");
        super.new(name);
    endfunction

    task body();
        super.body();
    endtask
endclass