typedef enum bit[7:0] {
    DUT_CHK   = 8'hCC
} dut_e;